module Seg(
	I,O
);

input [3:0]I;
output [6:0]O;

reg [6:0]O;

always @(1)
begin
	case(I)
			4'b0000:O=7'b1111110;
			4'b0001:O=7'b0110000;
			4'b0010:O=7'b1101101;
			4'b0011:O=7'b1111001;
			4'b0100:O=7'b0110011;
			4'b0101:O=7'b1011011;
			4'b0110:O=7'b1011111;
			4'b0111:O=7'b1110000;
			4'b1000:O=7'b1111111;
			4'b1001:O=7'b1110011;
			4'b1010:O=7'b1110111;
			4'b1011:O=7'b0011111;
			4'b1100:O=7'b1001110;
			4'b1101:O=7'b0111101;
			4'b1110:O=7'b1001111;
			4'b1111:O=7'b1000111;
			default:O=7'b0000000;  // Not in case
	endcase
end

endmodule
